//tb_data_buffer.sv

`timescale 1ns / 10ps

module tb_data_buffer();

  localparam CLK_PERIOD = 10;

  //DUT signals
  reg tb_clk;
  reg tb_n_rst;
  reg tb_clear;
  reg tb_store_rx_packet_data;
  reg [7:0] tb_rx_packet_data;
  reg tb_get_rx_data;
  reg [1:0] tb_data_size;
  reg [31:0] tb_tx_data;
  reg tb_store_tx_data;
  reg tb_get_tx_packet_data;
  reg tb_buffer_reserved;

  reg [6:0] tb_buffer_occupancy;
  reg [31:0] tb_rx_data;
  reg [7:0] tb_tx_packet_data;

  //*****************************************************************************
  // Clock Generation Block
  //*****************************************************************************
  // Clock generation block
  always begin
     // Start with clock low to avoid false rising edge events at t=0
     tb_clk = 1'b0;
     // Wait half of the clock period before toggling clock value (maintain 50% duty cycle)
     #(CLK_PERIOD/2.0);
     tb_clk = 1'b1;
     // Wait half of the clock period before toggling clock value via rerunning the block (maintain 50% duty cycle)
     #(CLK_PERIOD/2.0);
  end

  data_buffer DUT (.clk(tb_clk),
                   .n_rst(tb_n_rst),
                   .clear(tb_clear),
                   .store_rx_packet_data(tb_store_rx_packet_data),
                   .rx_packet_data(tb_rx_packet_data),
                   .get_rx_data(tb_get_rx_data),
                   .data_size(tb_data_size),
                   .tx_data(tb_tx_data),
                   .store_tx_data(tb_store_tx_data),
                   .get_tx_packet_data(tb_get_tx_packet_data),
                   .buffer_reserved(tb_buffer_reserved),
                   .buffer_occupancy(tb_buffer_occupancy),
                   .rx_data(tb_rx_data),
                   .tx_packet_data(tb_tx_packet_data));

   //*****************************************************************************
   // DUT Related TB Tasks
   //*****************************************************************************
   // Task for standard DUT reset procedure
   task reset_dut;
      begin
	 // Activate the reset
	 tb_n_rst = 1'b0;

	 // Maintain the reset for more than one cycle
	 @(posedge tb_clk);
	 @(posedge tb_clk);

	 // Wait until safely away from rising edge of the clock before releasing
	 @(negedge tb_clk);
	 tb_n_rst = 1'b1;

	 // Leave out of reset for a couple cycles before allowing other stimulus
	 // Wait for negative clock edges,
	 // since inputs to DUT should normally be applied away from rising clock edges
	 @(negedge tb_clk);
	 @(negedge tb_clk);
      end
   endtask // reset_dut

   //task for receiving a byte from RX
   task rx_send_byte;
      input logic [7:0] rx_byte;
      begin
	 tb_rx_packet_data = rx_byte;
	 tb_store_rx_packet_data = 1'b1;
	 
	 @(posedge tb_clk); //hold rx_packet_data high for one clock cycle

	 tb_store_rx_packet_data  = 1'b0;
      end   
   endtask // rx_send_byte

   //add task for sending multiple bytes to buffer
   task rx_send_bytes;
      input integer num_bytes;
      input logic [(num_bytes * 8 - 1):0] data;
      integer 				  i;
      integer 				  top_of_byte;
      
      begin
	 for (i = 0; i < num_bytes; i++)
	   begin
	      top_of_byte = ((i + 1) * 8) - 1;	      
	      rx_send_byte(data[top_of_byte: top_of_byte - 7]);
	   end
      end
   endtask // rx_send_bytes
   
   //task for sending data to AHB-Lite Slave
   task slave_request_data;
      input logic [1:0] data_size;
      input logic [31:0] expected_data;
      begin
	 tb_get_rx_data = 1'b1;
	 case(data_size)
	   2'd0: begin //1 byte
	      assert({24'd0, expected_data[7:0]} == tb_rx_data)
		$info("correct RX data for read 1 byte from data buffer");
	      else
		$error("correct RX data for read 1 byte from data buffer");
	   end
	   2'd1: begin //2 byte
	      assert({16'd0, expected_data[15:0]} == tb_rx_data)
		$info("correct RX data for read 2 bytes from data buffer");
	      else
		$error("correct RX data for read 2 bytes from data buffer");
	   end
	   2'd2: begin //3 byte
	      assert({8'd0, expected_data[23:0]} == tb_rx_data)
		$info("correct RX data for read 3 bytes from data buffer");
	      else
		$error("correct RX data for read 3 bytes from data buffer");
	   end
	   2'd3: begin //4 byte
	      assert(expected_data == tb_rx_data)
		$info("correct RX data for read 4 bytes from data buffer");
	      else
		$error("correct RX data for read 4 bytes from data buffer");
	   end
	 endcase // case (data_size)
      end
   endtask // slave_request_data 
	 
   //task for storing TX data
   task send_tx_data;
      input logic [1:0] num_bytes;
      input logic [31:0] tx_data;
      begin
	 tb_get_rx_data = 1'b1;
	 case(data_size)
	   2'd0: begin //1 byte
	      tb_store_tx_data = {24'd0, tx_data[7:0]};
	   end
	   2'd1: begin //2 byte
	      tb_store_tx_data = {16'd0, tx_data[15:0]};

	   end
	   2'd2: begin //3 byte
	      tb_store_tx_data = {8'd0, tx_data[23:0]};

	   end
	   2'd3: begin //4 byte
	      tb_store_tx_data = tx_data;
	   end
	 endcase // case (data_size)
      end
   endtask // send_tx_data
   
   //task for requesting TX data packet
   task request_tx_packet;
      input logic [7:0] expected_byte;
      begin
	 tb_get_tx_data_packet = 1'b1;
	 @(posedge tb_clk);//wait a clock cycle after asserting
	 assert(expected_byte == tb_tx_packet_data)
	   $info("correct tx_packet_data sent to usb tx");
	 else
	   $error("incorrect tx_packet_data sent to usb tx");
	 tb_get_tx_data_packet = 1'b0;
      end
   endtask
      
	 
   //task for checking buffer occupancy
   task check_buffer_occupancy;
      input logic [6:0] expected_occupancy;
      begin
	 assert(tb_buffer_occupancy == expected_occupancy)
	   $info("correct output for buffer occupancy");
	 else
	   $error("incorrect output for buffer occupancy");
      end
   endtask // check_buffer_occupancy
   
   //TODO add task for setting buffer reserved and trying to write
   
   //TODO write test cases and run tasks to check operation
   
 		
endmodule
